
module FIFO_Ctrl(
    input Clk,
    input Rst_n,
    input [10:0]ADC_Sample_Rate,    //������Ƶֵ�����������Ϊ1000KHz
    input ADC_Conv_Done,
    output reg Acq_Valid           //�ɼ���Ч��־
);
parameter NUMBER_SAMPLES = 1024;
reg Acq_Valid_r;    //�ɼ���Ч��־//Debug
reg [10:0]Acq_Div_Cnt;    //�ɼ���Ƶ������//Debug

//�������ʷ�Ƶ
always@(posedge Clk or negedge Rst_n)
begin
    if (!Rst_n)
        Acq_Div_Cnt <= 0;
    else if(Acq_Div_Cnt >= ADC_Sample_Rate)
        Acq_Div_Cnt <= 0;
    else if(ADC_Conv_Done)
        Acq_Div_Cnt <= Acq_Div_Cnt + 1;
    else
        Acq_Div_Cnt <= Acq_Div_Cnt;
end

//����������Ч��־,ֱ���ɼ����ݵ���Ŀ��ֵ���������ʶ
always@(posedge Clk or negedge Rst_n)
begin
    if (!Rst_n)
        Acq_Valid <= 0;
    else if(Acq_Div_Cnt >= ADC_Sample_Rate)
        Acq_Valid <= 1;
    else
        Acq_Valid <= 0;
end

endmodule