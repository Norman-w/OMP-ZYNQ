`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/07/27 16:48:31
// Design Name: 
// Module Name: AD7606_Driver
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module AD7606_Driver(
	Clk,
	Reset_n,
	Go,
	Speed_Set,
	Conv_Done,
	Channel_Set,
	ad7606_cs_n_o,   
	ad7606_rd_n_o,   
	ad7606_busy_i,   
	ad7606_db_i,     
	ad7606_os_o,     
	ad7606_reset_o,  
	ad7606_convst_o, 
	
	data_flag,
	data_mult_ch,
	ch_dat_valid
	
);

	input wire Clk;        //ʱ�ӣ�Ϊ���ò�������׼ȷ��Ҫ��Ϊ100MHz
	input wire Reset_n;    //��λ���͵�ƽ��λ
	input wire Go;         //����ʹ���źţ�Ϊ�ߵ�ƽ��ʹ�ܲ������͵�ƽ�����Ѿ���ʼ��һ�ֲ���������ֹͣ��һ�β�����
	input wire [25:0]Speed_Set; //�������ʿ��ƶ˿ڣ�Speed_Set = 100000000/speed - 1
	input wire [2:0]Channel_Set;//����ͨ�����ã��ɼ���0ͨ�����趨ͨ��Channel_Set��ֵ

	output reg Conv_Done;          //һ�β�����ɱ�־�źţ���ʱ�����������źš�ÿ��8��ͨ�����������󣬲���һ���������źš�

	output wire ad7606_cs_n_o;     //AD Ƭѡ�ź� ���Դ�AD7606�ж�ȡת�����ʱ����Ҫʹ���ź�Ϊ�͵�ƽ
	output reg ad7606_rd_n_o;      //AD �������ź�
	input wire ad7606_busy_i;      //AD æµ�ź�
	input wire [15:0]ad7606_db_i;  //AD �ɼ�������
	output wire [2:0]ad7606_os_o;  //AD OS����
	output reg ad7606_reset_o;     //AD ��λ�ź�
	output reg ad7606_convst_o;    //AD ת����ʼ�ź�
		
	/***
	��ͨ����������˿ڣ���ͨ��16λ���ڲ�ͬ��ʱ�̣������ͬͨ����ת�������ʹ��ʱ����data_flag�ź���ϣ�
    data_flag ����һλ���ָ����壬�����ǰdata_mult_ch��ֵΪ��ͨ����ת�������
    �ö˿���Ƶ�Ŀ����������FIFO��RAM �ȴ洢���д洢���ʱʹ�á�
	***/
	output reg [15:0]data_mult_ch;         //��ͨ����������˿�
	output reg [7:0]data_flag;             //8��ͨ����ת�������Ч��־�ź�
	
	output reg ch_dat_valid;

	assign ad7606_os_o = 0;                //��ʹ�ù�����
	assign ad7606_cs_n_o = ad7606_rd_n_o;  //���������ź����ӵ�Ƭѡ�ź�
	reg [7:0]state;                        //�������л�����
	reg [1:0]ad7606_busy_r;                //��¼busy�źŵ�ǰ������״̬
	
	//����ad7606_busy_r����λΪ�ϴ�ad7606_busy_i��״̬����λΪ����״̬
	always@(posedge Clk)
		ad7606_busy_r <= {ad7606_busy_r[0],ad7606_busy_i};
	
	//���������л��ļ���ֵ�õ���ǰ��Чͨ����־
	always@(posedge Clk or negedge Reset_n)
	if(!Reset_n)
		data_flag <= 0;
	else begin
		data_flag[0] <= state == 30;
		data_flag[1] <= state == 40;
		data_flag[2] <= state == 50;
		data_flag[3] <= state == 60;
		data_flag[4] <= state == 70;
		data_flag[5] <= state == 80;
		data_flag[6] <= state == 90;
		data_flag[7] <= state == 100;	
	end
	
	//��ÿ��ͨ�����ݲɼ���ɺ󣬽��µĲɼ�ֵ����
	always@(posedge Clk or negedge Reset_n)
	if(!Reset_n)
		data_mult_ch <= 0;
	else begin
		data_mult_ch <= 
			 (  (state == 30)
			 || (state == 40)
			 || (state == 50)
			 || (state == 60)
			 || (state == 70)
			 || (state == 80)
			 || (state == 90)
			 || (state == 100)
			)? ad7606_db_i:data_mult_ch;	
	end

	reg [25:0]cnt;     //������������cnt
	
	//����ֵÿ���ڼ�һ������������Speed_Setʱ������ֵ����
	always@(posedge Clk or negedge Reset_n)
	if(!Reset_n)
		cnt <= 0;
	else if(cnt == Speed_Set)
		cnt <= 0;
	else
		cnt <= cnt + 1'b1;
		
	wire trig = cnt == Speed_Set;  //��cnt=Speed_Setʱ��trig=1������Ϊ0
	
	//ʹ���������л�ģ��ʱ��ÿ�μ�����Speed_Setʱ��ȡ����
	always@(posedge Clk or negedge Reset_n)
	if(!Reset_n)begin
		state <= 0;
		ad7606_convst_o <= 1;
		Conv_Done <= 0;
		ad7606_rd_n_o <= 1;
		ad7606_reset_o <= 0;
	end
	else begin
		case(state)
			0:
				if(Go && trig)begin
					state <= 10;
					ad7606_convst_o <= 0;
					ad7606_rd_n_o <= 1;
					Conv_Done <= 0;
					ad7606_reset_o <= 0;
				end
				else begin
					state <= 0;
					ad7606_convst_o <= 1;
					ad7606_rd_n_o <= 1;
					ad7606_reset_o <= 0;
				end
					
			1: state <= state + 1'b1;
			2: state <= state + 1'b1;
			3: state <= state + 1'b1;
			4: state <= state + 1'b1;
			5: state <= state + 1'b1;
			6: state <= state + 1'b1;
			7: state <= state + 1'b1;
			8: state <= state + 1'b1;
			9: state <= state + 1'b1;
			10: state <= state + 1'b1;
			11: begin state <= state + 1'b1;ad7606_convst_o <= 1;end  //convst�����أ���������ת��
			12: begin state <= state + 1'b1;end
			13: state <= state + 1'b1;
			14: state <= state + 1'b1;
			15: state <= state + 1'b1;
			16: state <= state + 1'b1;
			17: state <= state + 1'b1;
			18: state <= state + 1'b1;
			19: if(ad7606_busy_r[1])state <= state;  //��ad7606_busy_i�ϴ�Ϊ��˵��ת��δ��ɣ���ѭ������״ֱ̬��ת�����
			    else begin state <= state + 3'd4;ad7606_rd_n_o <= 0;end  //���ϴ�ad7606_busy_iΪ�ͣ�˵����ת����ɣ����²������������14
			20: state <= state + 1'b1;
			21: state <= state + 1'b1;
			22: state <= state + 1'b1;
			23: state <= state + 1'b1;
			24: state <= state + 1'b1;
			25: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end
			26: state <= state + 1'b1;
			27: state <= state + 1'b1;
			28: state <= state + 1'b1;
			29: begin ad7606_rd_n_o <= 1; state <= state + 1'b1;end  // ad7606_rd_n_o�����أ����ɶ�ȡ��������
			30: state <= state + 1'b1;
			31: state <= state + 1'b1;
			32: state <= state + 1'b1;
			33: state <= state + 1'b1;
			34: state <= state + 1'b1;
			35: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			36: begin state <= state + 1'b1;end  
			37: begin state <= state + 1'b1;end
			38: begin state <= state + 1'b1;end
			39: begin ad7606_rd_n_o <= 1; state <= state + 1'b1;end  //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			40: state <= state + 1'b1;
			41: state <= state + 1'b1;
			42: state <= state + 1'b1;
			43: state <= state + 1'b1;
			44: state <= state + 1'b1;
			45: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			46: state <= state + 1'b1;
			47: begin state <= state + 1'b1;end
			48: begin state <= state + 1'b1;end
			49: begin ad7606_rd_n_o <= 1;  state <= state + 1'b1;end //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			50: state <= state + 1'b1;
			51: state <= state + 1'b1;
			52: state <= state + 1'b1;
			53: state <= state + 1'b1;
			54: state <= state + 1'b1;
			55: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			56: state <= state + 1'b1;
			57: begin state <= state + 1'b1;end
			58: begin state <= state + 1'b1;end
			59: begin ad7606_rd_n_o <= 1;  state <= state + 1'b1;end //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			60: state <= state + 1'b1;
			61: state <= state + 1'b1;
			62: state <= state + 1'b1;
			63: state <= state + 1'b1;
			64: state <= state + 1'b1;
			65: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			66: state <= state + 1'b1;
			67: begin state <= state + 1'b1;end
			68: begin state <= state + 1'b1;end
			69: begin ad7606_rd_n_o <= 1;  state <= state + 1'b1;end //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			70: state <= state + 1'b1;
			71: state <= state + 1'b1;
			72: state <= state + 1'b1;
			73: state <= state + 1'b1;
			74: state <= state + 1'b1;
			75: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			76: state <= state + 1'b1;
			77: begin state <= state + 1'b1;end
			78: begin state <= state + 1'b1;end
			79: begin ad7606_rd_n_o <= 1;  state <= state + 1'b1;end //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			80: state <= state + 1'b1;
			81: state <= state + 1'b1;
			82: state <= state + 1'b1;
			83: state <= state + 1'b1;
			84: state <= state + 1'b1;
			85: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			86: state <= state + 1'b1;
			87: begin state <= state + 1'b1;end
			88: begin state <= state + 1'b1;end
			89: begin ad7606_rd_n_o <= 1; state <= state + 1'b1;end //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			90: state <= state + 1'b1;
			91: state <= state + 1'b1;
			92: state <= state + 1'b1;
			93: state <= state + 1'b1;
			94: state <= state + 1'b1;
			95: begin ad7606_rd_n_o <= 0; state <= state + 1'b1;end  //ad7606_rd_n_o�½��أ����²������
			96: state <= state + 1'b1;
			97: begin state <= state + 1'b1;end
			98: begin state <= state + 1'b1;end
			99: begin ad7606_rd_n_o <= 1;  state <= state + 1'b1;end //ad7606_rd_n_o�����أ����ɶ�ȡ��������
			100: begin state <= state + 1'b1; Conv_Done <= 1; end    //ת������ź�Conv_Done��Ϊ�ߵ�ƽ
			101: begin state <= state + 1'b1; ad7606_reset_o <= 1; Conv_Done <= 0; end//��λad7606�ڲ��������ܵ�Ԫ�Ĺ���״̬,Conv_Done��Ϊ�͵�ƽ
			102: begin state <= 0;ad7606_reset_o <= 0; end    //ad7606_reset_o��ߣ�state����
			default:
				begin
					state <= 0;
					ad7606_convst_o <= 1;
					Conv_Done <= 0;
					ad7606_rd_n_o <= 1;
					ad7606_reset_o <= 0;
				end
		endcase
	end
	
	//���������л��ļ���ֵ�õ�stream��������ź�
	always@(posedge Clk or negedge Reset_n)
	if(!Reset_n)
		ch_dat_valid <= 0;
	else if(state==(Channel_Set+3)*10)
        ch_dat_valid <= 1;
	else
        ch_dat_valid <= 0;
        
    

endmodule


