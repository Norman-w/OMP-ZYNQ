`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/11/29 18:22:24
// Design Name: 
// Module Name: ADC_Measure_Freq
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: ����ADC��������ĵ�ѹƵ��
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ADC_Measure_Freq(
    input Clk,
    input Rst_n,
    input signed [15:0]Trig_Val,       //����ֵ
    input signed [15:0]ADC_Data,       //ADC����
    input ADC_Conv_Done,        //ADC���βɼ�����ź�
    output reg [31:0]Freq_Val  //Ƶ�ʲ���ֵ
);
parameter TIME_CNT_VAL = 99999999; //�趨����ֵ�����Ʋ���ʱ��
reg signed [15:0]ADC_Data_Pre;   //������һ������ֵ
reg ADC_Conv_Done_r;      //���βɼ�����źŴ���
reg [31:0]Time_Cnt;       //ʱ�������
reg [31:0]Cycle_Cnt_Pre;  //������һ������ֵ
reg signed [15:0]Trig_Val_r;     //�洢����ֵ����ֹ��;�ı�
reg [31:0]Cycle_Cnt; //���ڼ�����
reg [31:0]Freq_Add;   //��λʱ����Ƶ���ۼ�

//����1��
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        Time_Cnt <= 0;
    else if(Time_Cnt >= TIME_CNT_VAL)
		Time_Cnt <= 0;
    else
        Time_Cnt <= Time_Cnt + 1;
end

//1�����ۼӴ����������Դ˲��Ƶ��
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        Freq_Add <= 0;
	else if(Time_Cnt >= TIME_CNT_VAL)
		Freq_Add <= 0;
	else if((ADC_Data_Pre <= Trig_Val_r) && (ADC_Data >= Trig_Val_r) && (ADC_Data_Pre < ADC_Data) && ADC_Conv_Done) begin
        if(Cycle_Cnt <= Cycle_Cnt_Pre[31:1])//��ǰ���ڼ���С�ڵ�����һ���������ڵ�һ�룬��˴δ����쳣������������Ч
            Freq_Add <= Freq_Add;
        else 
            Freq_Add <= Freq_Add + 1;
    end
	else
        Freq_Add <= Freq_Add;
end

//��¼һ�δ������ڵ�ʱ��
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        Cycle_Cnt <= 0;
    else if((ADC_Data_Pre <= Trig_Val_r) && (ADC_Data >= Trig_Val_r) && (ADC_Data_Pre < ADC_Data) && ADC_Conv_Done)
		Cycle_Cnt <= 0;
    else
        Cycle_Cnt <= Cycle_Cnt + 1;
end

//������һ�δ������ڵ�ʱ��
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        Cycle_Cnt_Pre <= 0;
    else if((ADC_Data_Pre <= Trig_Val_r) && (ADC_Data >= Trig_Val_r) && (ADC_Data_Pre < ADC_Data) && ADC_Conv_Done)
		Cycle_Cnt_Pre <= Cycle_Cnt;
    else
        Cycle_Cnt_Pre <= Cycle_Cnt_Pre;
end

//���津���趨ֵ����ֹ��;���޸ģ�ÿ�β���һ���������޸�
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        Trig_Val_r <= 0;
    else if(Time_Cnt >= TIME_CNT_VAL)
		Trig_Val_r <= Trig_Val;
    else
        Trig_Val_r <= Trig_Val_r;
end

//������һ��ADC����ֵ
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n) begin
        ADC_Data_Pre <= 0;
    end
    else if(ADC_Conv_Done) begin
        ADC_Data_Pre <= ADC_Data;
    end
    else begin
        ADC_Data_Pre <= ADC_Data_Pre;
    end
end

//ADC����ת������źŴ���
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        ADC_Conv_Done_r <= 0;
    else
        ADC_Conv_Done_r <= ADC_Conv_Done;
end

//����1����������Ƶ��
always@(posedge Clk or negedge Rst_n)
begin
    if(!Rst_n)
        Freq_Val <= 0;
	else if(Time_Cnt >= TIME_CNT_VAL)
	    Freq_Val <= Freq_Add;
    else
        Freq_Val <= Freq_Val;
end

endmodule
