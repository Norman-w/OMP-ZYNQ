`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/11/29 18:22:24
// Design Name: 
// Module Name: ADC128S102
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ADC128S102(
			Clk,
			Rst_n,
			
			Channel,
			Data,
			
			En_Conv,
			Conv_Done,
			ADC_State,
			DIV_PARAM,
			
			ADC_SCLK,
			ADC_DOUT,
			ADC_DIN,
			ADC_CS_N	
		);

	input Clk;	//����ʱ��
	input Rst_n; //��λ���룬�͵�ƽ��λ
	input [2:0]Channel;	//ADCת��ͨ��ѡ��
	output reg [11:0]Data;	//ADCת�����
	
	input En_Conv;	//ʹ�ܵ���ת�������ź�Ϊ��������Ч��������ʹ��һ��ת��
	output reg Conv_Done;	//ת������źţ����ת�������һ��ʱ�����ڵĸ�����
	output ADC_State;	//ADC����״̬��ADC����ת��ʱΪ�͵�ƽ������ʱΪ�ߵ�ƽ
	input [7:0]DIV_PARAM;	//ʱ�ӷ�Ƶ���ã�ʵ��SCLKʱ�� Ƶ�� = fclk / ��DIV_PARAM * 2��
	
	output reg ADC_SCLK;	//ADC �������ݽӿ�ʱ���ź�
	output reg ADC_CS_N;  //ADC �������ݽӿ�ʹ���ź�
	input  ADC_DOUT;		//ADCת���������ADC���FPGA
	output reg ADC_DIN;	//ADC�����ź��������FPGA����ͨ�������ָ�ADC
	
	reg [2:0]r_Channel; //ͨ��ѡ���ڲ��Ĵ���
	reg [11:0]r_data;	//ת�������ȡ�ڲ��Ĵ���
	
	reg [7:0]DIV_CNT;//��Ƶ������
	reg SCLK2X;//2��SCLK�Ĳ���ʱ��
	
	reg [5:0]SCLK_GEN_CNT;//SCLK���������л�������

	
	reg en;//ת��ʹ���ź�
	
	//��ÿ��ʹ��ת����ʱ�򣬼Ĵ�Channel��ֵ����ֹ��ת�������и�ֵ�����仯
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		r_Channel <= 3'd0;
	else if(En_Conv)
		r_Channel <= Channel;
	else
		r_Channel <= r_Channel;

	//����ʹ��ת���ź�
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		en  <= 1'b0;
	else if(En_Conv)
		en  <= 1'b1;
	else if(Conv_Done)
		en  <= 1'b0;
	else
		en  <= en;
		
	//����2��SCLKʹ��ʱ�Ӽ�����
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		DIV_CNT  <= 8'd0;
	else if(en)begin
		if(DIV_CNT >= (DIV_PARAM - 1'b1))
			DIV_CNT  <= 8'd0;
		else 
			DIV_CNT  <= DIV_CNT + 1'b1;
	end else	
		DIV_CNT  <= 8'd0;

	//����2��SCLKʹ��ʱ��
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		SCLK2X  <= 1'b0;
	else if(en && (DIV_CNT >= (DIV_PARAM - 1'b1)))
		SCLK2X  <= 1'b1;
	else
		SCLK2X  <= 1'b0;
		
	//�������м�����
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)
		SCLK_GEN_CNT  <= 6'd0;
	else if(SCLK2X && en)begin
		if(SCLK_GEN_CNT >= 6'd31)
			SCLK_GEN_CNT  <= 6'd0;
		else
			SCLK_GEN_CNT  <= SCLK_GEN_CNT + 1'd1;
	end else
		SCLK_GEN_CNT  <= SCLK_GEN_CNT;
	
	//���л�ʵ��ADC�������ݽӿڵ����ݷ��ͺͽ���	
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)begin
		ADC_SCLK <= 1'b1;
		ADC_CS_N <= 1'b1;
		ADC_DIN  <= 1'b1;
	end else if(en) begin
		if(SCLK2X)begin
			case(SCLK_GEN_CNT)
				6'd0:begin ADC_SCLK <= 1'b0; ADC_DIN  <= 1'b0; end
				6'd1:begin ADC_SCLK <= 1'b1; end
				6'd2:begin ADC_SCLK <= 1'b0; end
				6'd3:begin ADC_SCLK <= 1'b1; end
				6'd4:begin ADC_SCLK <= 1'b0; ADC_DIN  <= r_Channel[2];end	//addr[2]
				6'd5:begin ADC_SCLK <= 1'b1; end
				6'd6:begin ADC_SCLK <= 1'b0; ADC_DIN  <= r_Channel[1];end	//addr[1]
				6'd7:begin ADC_SCLK <= 1'b1; end
				6'd8:begin ADC_SCLK <= 1'b0; ADC_DIN  <= r_Channel[0];end	//addr[0]

				//ÿ�������أ��Ĵ�ADC��������������ϵ�ת�����
				6'd9,6'd11,6'd13,6'd15,6'd17,6'd19,6'd21,6'd23,6'd25,6'd27,6'd29,6'd31:
					begin ADC_SCLK <= 1'b1; r_data <= {r_data[10:0], ADC_DOUT}; end	//ѭ����λ�Ĵ�DOUT�ϵ�12������
				
				6'd10,6'd12,6'd14,6'd16,6'd18,6'd20,6'd22,6'd24,6'd26,6'd28,6'd30:
					begin ADC_SCLK <= 1'b0; end

				default:begin ADC_CS_N <= 1'b0; end //��ת��������
			endcase
		end
		else ;
	end else begin
		ADC_CS_N <= 1'b0;
	end
	
	//ת�����ʱ����ת����������Data�˿ڣ�ͬʱ����һ��ʱ�����ڵĸ������ź�
	always@(posedge Clk or negedge Rst_n)
	if(!Rst_n)begin
		Data <= 12'd0; 
		Conv_Done <= 1'b0;
	end else if(en && (SCLK2X == 1'b1) && (SCLK_GEN_CNT >= 6'd31))begin
		Data <= {r_data[10:0], ADC_DOUT}; 
		Conv_Done <= 1'b1;
	end else begin
		Data <= Data; 
		Conv_Done <= 1'b0;
	end
	
	//����ADC����״ָ̬ʾ�ź�
	assign ADC_State = ADC_CS_N;

endmodule
